module CNN (
input [2:0] x,
output [0:0] y
);
endmodule
