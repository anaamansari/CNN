module input_configure # (

I= 32,
O= 32,

N=32,
Q=15,

L1=4,L2=24,L3=6,L4=6,L5=16 
)

(
input [N-1:0] IN [I-1:0],
output [N-1:0] OUT [O-1:0]
);



endmodule 