module PE_cont
(
	input Tn,
	input Tm,
	
	output Benes_config,
	output PE_enable

);

endmodule
